
module block_move (iCLK, reset, in, out);
